`include "classa.sv"
class B;

    A obj_a=new;
    function new(); 
    obj_a.print(5);
    A::print(10);
    endfunction
    
endclass:B


