`include "classb.sv"
module example;
  B obj_b;  
  initial begin
    obj_b = new();
  end
endmodule
